module direct_cache #(parameter LINE_LENGTH, CACHE_LENGTH, ADDRESS_SIZE)();

endmodule
